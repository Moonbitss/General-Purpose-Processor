library verilog;
use verilog.vl_types.all;
entity ALU2basic_vlg_vec_tst is
end ALU2basic_vlg_vec_tst;
