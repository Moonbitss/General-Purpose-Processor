library verilog;
use verilog.vl_types.all;
entity ALU2Block_vlg_vec_tst is
end ALU2Block_vlg_vec_tst;
