library verilog;
use verilog.vl_types.all;
entity ALU3block_vlg_vec_tst is
end ALU3block_vlg_vec_tst;
