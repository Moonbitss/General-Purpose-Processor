library verilog;
use verilog.vl_types.all;
entity Part1ALU_vlg_vec_tst is
end Part1ALU_vlg_vec_tst;
