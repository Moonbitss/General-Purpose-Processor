library verilog;
use verilog.vl_types.all;
entity decode4to16_vlg_vec_tst is
end decode4to16_vlg_vec_tst;
