library verilog;
use verilog.vl_types.all;
entity ALUbasic_vlg_vec_tst is
end ALUbasic_vlg_vec_tst;
