library verilog;
use verilog.vl_types.all;
entity ssegblock_vlg_vec_tst is
end ssegblock_vlg_vec_tst;
